<?xml version="1.0" encoding="UTF-8"?><Batch version="2.0"><TaskList><Task type="ResizeCanvasByAspectRatioTask" enabled="true"><AspectRatio>1:1</AspectRatio><Justification>4</Justification><MainSide>1</MainSide><BackColor>#FFFFFF</BackColor><FillType>0</FillType><Alpha>255</Alpha></Task><Task type="ResizeTask" enabled="true"><Width units="0"><![CDATA[5120]]></Width><Height units="0"><![CDATA[5120]]></Height><DPI><![CDATA[-1]]></DPI><Filter>9</Filter><UseProportions>False</UseProportions><ResizeType>0</ResizeType><ProportionsSize>0</ProportionsSize></Task><Task type="RoundImageTask" enabled="true"><RoundWidth units="0">1000</RoundWidth><RoundHeight units="0">1000</RoundHeight><RoundBackground>#000000</RoundBackground><RoundBackTransp>-1</RoundBackTransp></Task><Task type="ResizeTask" enabled="true"><Width units="0"><![CDATA[256]]></Width><Height units="0"><![CDATA[256]]></Height><DPI><![CDATA[-1]]></DPI><Filter>9</Filter><UseProportions>True</UseProportions><ResizeType>0</ResizeType><ProportionsSize>0</ProportionsSize></Task><Task type="SaveAsTask" enabled="true"><FileName><![CDATA[<Original Name (Without Extension)>]]></FileName><PreserveStruct>False</PreserveStruct><CommonFolder><![CDATA[]]></CommonFolder><FileType>PNG</FileType><FilePath><![CDATA[C:\Users\thomt\AppData\Roaming\Tapstream\icons]]></FilePath><FileExists>0</FileExists><DefaultOptions>True</DefaultOptions><BMPCompression>0</BMPCompression><BMPVersion>1</BMPVersion><JPEGColorSpace>2</JPEGColorSpace><JPEGDCTMethod>0</JPEGDCTMethod><JPEGCromaSubsampling>1</JPEGCromaSubsampling><JPEGOptimalHuffman>False</JPEGOptimalHuffman><JPEGQuality>95</JPEGQuality><PNGCompression>5</PNGCompression><PNGFilter>1</PNGFilter><PNGInterlaced>False</PNGInterlaced><J2000ColorSpace>1</J2000ColorSpace><J2000Rate>0.500</J2000Rate><PCXCompression>1</PCXCompression><HDPLossless>False</HDPLossless><HDPImageQuality>0.900</HDPImageQuality><TGACompressed>False</TGACompressed><DDSMIPLevels>8</DDSMIPLevels><DDSMipMapFilter>4</DDSMipMapFilter><DDSFormat>71</DDSFormat><TIFFCompression>0</TIFFCompression><TIFFJPEGColorSpace>2</TIFFJPEGColorSpace><TIFFJPEGQuality>95</TIFFJPEGQuality><TIFFZIPCompression>1</TIFFZIPCompression><TIFFPlanarConf>1</TIFFPlanarConf><DICOMCompression>6</DICOMCompression><DICOMJPEG2000Rate>1</DICOMJPEG2000Rate><DICOMJPEGQuality>95</DICOMJPEGQuality><WEBPLossless>0</WEBPLossless><WEBPQuality>75</WEBPQuality><WEBPMethod>0</WEBPMethod><WEBPTargetSize>0</WEBPTargetSize><WEBPFilterStrength>0</WEBPFilterStrength><WEBPFilterSharpness>0</WEBPFilterSharpness></Task></TaskList></Batch>